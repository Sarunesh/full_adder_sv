mailbox gen2bfm = new();
mailbox mon2cov = new();
mailbox mon2sbd = new();
