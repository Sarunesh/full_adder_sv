`include "fa_common.sv"
`include "fa_tx.sv"
`include "full_adder.v"
`include "fa_interface.sv"
`include "fa_bfm.sv"
`include "fa_cov.sv"
`include "fa_gen.sv"
`include "fa_mon.sv"
`include "fa_sbd.sv"
`include "fa_agent.sv"
`include "fa_env.sv"
`include "top.sv"
