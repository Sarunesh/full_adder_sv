mailbox gen2bfm = new();
mailbox mon2cov = new();
mailbox mon2sbd = new();

class fa_common;
	static int count=30;
	static int bfm_count;
	static int gen_count;
  	static int sum_match;
	static int sum_mismatch;
	static int carry_match;
	static int carry_mismatch;
endclass
